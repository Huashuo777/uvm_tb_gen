adsad

dfadf
dfaf
