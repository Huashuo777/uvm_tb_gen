ddddddddddddddadsad

dfadf
dfaf
