//----------------------------------------------------------------------------------
// This code is copyrighted by BrentWang and cannot be used for commercial purposes
// The github address:https://github.com/brentwang-lab/uvm_tb_gen                   
// You can refer to the book <UVM Experiment Guide> for learning, this is on this github
// If you have any questions, please contact email:brent_wang@foxmail.com          
//----------------------------------------------------------------------------------
//                                                                                  
// Author  : BrentWang                                                              
// Project : UVM study                                                              
// Date    : Sat Jan 26 06:05:52 WAT 2022                                           
//----------------------------------------------------------------------------------
//                                                                                  
// Description:                                                                     
//     File for apb_env_pkg.sv                                                       
//----------------------------------------------------------------------------------
`ifndef APB_ENV_PKG__SV
`define APB_ENV_PKG__SV
`include "apb_define.sv"
`include "apb_env_interface.sv"
package apb_env_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "apb_common_include.svh"
    `include "apb_master_include.svh"
    `include "apb_slave_include.svh"
    `include "apb_env_config.sv"
    `include "apb_virtual_sequencer.sv"
    `include "apb_virtual_sequence.sv"
    `include "apb_environment.sv"
endpackage : apb_env_pkg
`endif //APB_ENV_PKG__SV
