//----------------------------------------------------------------------------------
// This code is copyrighted by BrentWang and cannot be used for commercial purposes
// The github address:https://github.com/brentwang-lab/uvm_tb_gen                   
// You can refer to the book <UVM Experiment Guide> for learning, this is on this github
// If you have any questions, please contact email:brent_wang@foxmail.com          
//----------------------------------------------------------------------------------
//                                                                                  
// Author  : BrentWang                                                              
// Project : UVM study                                                              
// Date    : Sat Jan 26 06:05:52 WAT 2022                                           
//----------------------------------------------------------------------------------
//                                                                                  
// Description:                                                                     
//     File for apb_common_include.svh                                                       
//----------------------------------------------------------------------------------
`ifndef APB_COMMON_INCLUDE__SV
`define APB_COMMON_INCLUDE__SV
    `include "apb_type.sv"
    `include "apb_base_config.sv"
    `include "apb_base_item.sv" 
`endif //APB_COMMON_INCLUDE__SV
