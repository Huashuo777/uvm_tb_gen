//----------------------------------------------------------------------------------
// This code is copyrighted by BrentWang and cannot be used for commercial purposes
// The github address:https://github.com/brentwang-lab/uvm_tb_gen                   
// You can refer to the book <UVM Experiment Guide> for learning, this is on this github
// If you have any questions, please contact email:brent_wang@foxmail.com          
//----------------------------------------------------------------------------------
//                                                                                  
// Author  : BrentWang                                                              
// Project : UVM study                                                              
// Date    : Sat Jan 26 06:05:52 WAT 2022                                           
//----------------------------------------------------------------------------------
//                                                                                  
// Description:                                                                     
//     File for dadd_include.svh                                                       
//----------------------------------------------------------------------------------
`include "dadd_item.sv"
`include "dadd_driver.sv"
`include "dadd_imonitor.sv"
`include "dadd_sequencer.sv"
`include "dadd_iagent.sv"
`include "dadd_omonitor.sv"
`include "dadd_oagent.sv"
