//----------------------------------------------------------------------------------
// This code is copyrighted by BrentWang and cannot be used for commercial purposes
// The github address:https://github.com/brentwang-lab/uvm_tb_gen                   
// You can refer to the book <UVM Experiment Guide> for learning, this is on this github
// If you have any questions, please contact email:brent_wang@foxmail.com          
//----------------------------------------------------------------------------------
//                                                                                  
// Author  : BrentWang                                                              
// Project : UVM study                                                              
// Date    : Sat Jan 26 06:05:52 WAT 2022                                           
//----------------------------------------------------------------------------------
//                                                                                  
// Description:                                                                     
//     File for dadd_loc_include.svh                                                       
//----------------------------------------------------------------------------------
`ifndef DADD_LOC_INCLUDE__SVH
`define DADD_LOC_INCLUDE__SVH
    `include "dadd_loc_item.sv"
    `include "dadd_loc_sequencer.sv"
    `include "dadd_loc_base_sequence.sv"
    `include "dadd_loc_driver.sv"
    `include "dadd_loc_imonitor.sv"
    `include "dadd_loc_iagent.sv"
    `include "dadd_loc_omonitor.sv"
    `include "dadd_loc_oagent.sv"
`endif // DADD_LOC_INCLUDE__SVH
